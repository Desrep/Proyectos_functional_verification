`include "interface.sv"
`include "stimulus.sv"
`include "scoreboard.sv"
`include "driver.sv"
`include "monitor.sv"
`include "coverage.sv"
`include "env.sv"
//`include "test1.sv"
`include "test2.sv"
`include "top.sv"
`include "assertions.sv"

