
`include "interface.sv"
`include "seq_item.sv"
`include "sequencer.sv"
`include "sequence.sv"
`include "driver.sv"
`include "monitor.sv"
`include "monitor_decode.sv"
`include "monitor_decode_column.sv"
`include "agent.sv"
`include "agent_passive.sv"
`include "agent_passive_col.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "test.sv"
`include "wr_rd_test.sv"
`include "tb_top.sv"
`include "coverage.sv"


